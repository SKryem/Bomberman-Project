// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen Apr  2023  
// (c) Technion IIT, Department of Electrical Engineering 2023 



module	explosionMineMatrixBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic OneSecPulse,
					input logic mineExploded,
					
					
					
					output logic [3:0] explosionIndexX,
					output logic [3:0] explosionIndexY,
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap

 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */

// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 16*16 and use only the top left 16*15 squares 
// this is the bitmap  of the maze , if there is a specific value  the  whole 32*32 rectange will be drawn on the screen
// there are  16 options of differents kinds of 32*32 squares 
// all numbers here are hard coded to simplify the  understanding 




const logic [0:15] [0:15] [3:0]  initial_map = {
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},// last line in home screen
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00}};
logic [0:15] [0:15] [3:0]  mineBitMapMask_p = initial_map;
logic [0:15] [0:15] [3:0]  mineBitMapMask_n;  

logic[0:31][0:31][7:0] object_colors = {
	{8'hda,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hda,8'hb6,8'hb6,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hb6,8'hb6,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hba},
	{8'hb6,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h25,8'h25,8'h25,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hda},
	{8'hb6,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'hda,8'h25,8'h25,8'h25,8'h25,8'h25,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hda},
	{8'hda,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h25,8'h24,8'hda,8'h6d,8'h25,8'h25,8'h25,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hda},
	{8'hda,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h25,8'h25,8'hda,8'h6d,8'h24,8'h25,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hda},
	{8'hb6,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h25,8'h25,8'h25,8'h25,8'h25,8'hb6,8'h24,8'h24,8'h65,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hda},
	{8'hb6,8'h24,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h24,8'h25,8'h25,8'h25,8'h25,8'h25,8'h91,8'hda,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hda,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hda},
	{8'hb6,8'h24,8'h24,8'h24,8'h24,8'h24,8'h6d,8'hb6,8'h91,8'h25,8'h24,8'h25,8'h25,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h25,8'h2d,8'h91,8'hb6,8'h91,8'h2c,8'h25,8'h6d,8'h6d,8'h6d,8'h6d,8'hda},
	{8'hba,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h91,8'hb6,8'h6d,8'h24,8'h6d,8'h6d,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h25,8'h24,8'hda,8'h91,8'h6d,8'h25,8'h25,8'h6d,8'h6d,8'h6d,8'h6d,8'hda},
	{8'hba,8'h24,8'h24,8'h24,8'h25,8'h25,8'h25,8'h25,8'h6d,8'h91,8'h91,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hda},
	{8'hba,8'h24,8'h24,8'h25,8'h25,8'h25,8'h25,8'h25,8'h24,8'h91,8'hda,8'h91,8'hb6,8'hb6,8'h91,8'hb6,8'h91,8'h91,8'h6d,8'h6d,8'hda,8'h91,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h2d,8'hda},
	{8'hda,8'h24,8'h25,8'h25,8'h25,8'h25,8'h25,8'h65,8'h6d,8'hb6,8'h6d,8'hff,8'h91,8'h6d,8'hb6,8'hb6,8'hb6,8'h91,8'h6d,8'hda,8'h6d,8'h6d,8'h6d,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h2d,8'h25,8'hda},
	{8'hda,8'h24,8'h25,8'h25,8'h25,8'h25,8'h6d,8'h6d,8'h6d,8'hb6,8'hb6,8'h91,8'hda,8'h6d,8'hb6,8'h91,8'hb6,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h25,8'h6d,8'h6d,8'h6d,8'h25,8'h25,8'h25,8'hda},
	{8'hda,8'h25,8'h25,8'h25,8'h25,8'h6d,8'h6d,8'h6d,8'h91,8'hb6,8'hb6,8'h6d,8'h6d,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6c,8'h24,8'h6d,8'h6d,8'h25,8'h25,8'h25,8'h25,8'hda},
	{8'hda,8'h25,8'h25,8'h25,8'h6d,8'h6d,8'hda,8'h6d,8'h91,8'hb6,8'h91,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h6d,8'h6d,8'h91,8'h6d,8'h6d,8'h24,8'hda,8'h25,8'h25,8'h25,8'h24,8'h25,8'hda},
	{8'hda,8'h25,8'hb6,8'hda,8'hda,8'hb6,8'hda,8'h6d,8'h6d,8'h91,8'hb6,8'hb6,8'h91,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'hda,8'hb6,8'hda,8'hda,8'h24,8'h25,8'hda},
	{8'hda,8'h25,8'h6d,8'h6d,8'h6d,8'h24,8'h91,8'h6d,8'h6d,8'h91,8'h91,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h91,8'h25,8'h6d,8'h6d,8'h6d,8'h25,8'hda},
	{8'hda,8'h2d,8'h6d,8'h6d,8'h25,8'h25,8'h6d,8'h6d,8'h6d,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h91,8'h6d,8'h6d,8'h24,8'h24,8'h6d,8'h20,8'h24,8'h24,8'h24,8'h24,8'hda},
	{8'hda,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h6d,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h25,8'h25,8'h25,8'h25,8'hda},
	{8'hda,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h65,8'h6d,8'h6d,8'h6d,8'hff,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'hda,8'h24,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h25,8'h25,8'h25,8'h25,8'h25,8'hda},
	{8'hda,8'h6d,8'h6d,8'h6d,8'h6d,8'h65,8'h25,8'h25,8'h6d,8'h6d,8'hda,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h91,8'h24,8'h24,8'hff,8'h24,8'h24,8'h24,8'h24,8'h25,8'h25,8'h25,8'h25,8'h25,8'h24,8'hda},
	{8'hda,8'h6d,8'h6d,8'h65,8'h25,8'h25,8'h25,8'h24,8'h24,8'h24,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h6d,8'h24,8'h24,8'hff,8'h24,8'h24,8'h24,8'h25,8'h25,8'h25,8'h24,8'h24,8'h24,8'hda},
	{8'hb6,8'h6d,8'h65,8'h25,8'h25,8'h25,8'h25,8'h71,8'hda,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h24,8'h25,8'h25,8'h24,8'h24,8'h24,8'h24,8'hda},
	{8'hb6,8'h65,8'h25,8'h25,8'h25,8'h25,8'h25,8'hb6,8'h91,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h25,8'h24,8'h24,8'h24,8'h24,8'h24,8'hda},
	{8'hb6,8'h25,8'h25,8'h25,8'h25,8'h24,8'hda,8'h6d,8'h25,8'h20,8'h24,8'h25,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'hda},
	{8'hb6,8'h25,8'h25,8'h25,8'h25,8'h24,8'h91,8'h6d,8'h24,8'h25,8'h25,8'h24,8'h25,8'h25,8'hdb,8'h91,8'h91,8'h6d,8'h24,8'h24,8'h25,8'h25,8'h25,8'h25,8'h6d,8'h6d,8'h00,8'h24,8'h24,8'h24,8'h20,8'hda},
	{8'hb6,8'h25,8'h25,8'h25,8'h25,8'h25,8'h24,8'h24,8'h24,8'h25,8'h25,8'h25,8'h25,8'h25,8'h24,8'h6d,8'h24,8'h24,8'h24,8'h25,8'h25,8'h25,8'h25,8'h24,8'h24,8'h00,8'h00,8'h24,8'h24,8'h24,8'h20,8'hda},
	{8'hb6,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h91,8'h6d,8'h24,8'h25,8'h25,8'h25,8'h25,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h20,8'hda},
	{8'hb6,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h6d,8'h6d,8'h24,8'h25,8'h25,8'h25,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h20,8'hda},
	{8'hb6,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h6d,8'h24,8'h25,8'h25,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h20,8'hda},
	{8'hda,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'hda},
	{8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hb6}};

 // pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <= TRANSPARENT_ENCODING ;
		mineBitMapMask_p = initial_map;

	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 
		mineBitMapMask_p <= mineBitMapMask_n;

		if ((InsideRectangle == 1'b1 )		& 	// only if inside the external bracket 
		   (mineBitMapMask_p[offsetY[8:5] ][offsetX[8:5]] > 4'h0 ))begin
						// take bits 5,6,7,8,9,10 from address to select  position in the maze    
						RGBout <= object_colors[offsetY[4:0]][offsetX[4:0]] ; 
		end
	end	
end

always_comb begin 

	mineBitMapMask_n = mineBitMapMask_p;
	
	if(mineExploded) begin
		mineBitMapMask_n[offsetY[8:5] ][offsetX[8:5]] = 0; // remove mine
	end
	
end


//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign explosionIndexX = offsetX[8:5];
assign explosionIndexY = offsetY[8:5];
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule

