// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen Apr  2023  
// (c) Technion IIT, Department of Electrical Engineering 2023 



module	explosionMatrixBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
		
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic [3:0] bombExplosionIndexX,
					input logic [3:0] bombExplosionIndexY,
					input logic [3:0] landMineExplosionIndexX,
					input logic [3:0] landMineExplosionIndexY,
					input logic [3:0] explosionMineExplosionIndexX,
					input logic [3:0] explosionMineExplosionIndexY,
					
					input logic explodeBomb,
					input logic random_dir, // random direction for explosion, 0 for vertical and 1 for horizontal
					input logic mineTriggered,// when the character steps on a mine
					input logic mineExploded, // when a bomb detonates a mine
					input logic OneSecPulse, 
					
					// output for explosion, 
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;
 
 
logic last_direction_p; // save last 4 explosions directions
logic last_direction_n;


// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */


// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 16*16 and use only the top left 16*15 squares 
// this is the bitmap  of the maze , if there is a specific value  the  whole 32*32 rectange will be drawn on the screen
// there are  16 options of differents kinds of 32*32 squares 
// all numbers here are hard coded to simplify the  understanding 


// start the bit map with zeroes, each value represents the timer remaining for the bomb to explode, 0-> no bomb



	const int explosion_length = 2;
	logic bombExplosion_executed_p;
	logic bombExplosion_executed_n;
	logic landMineExplosion_executed_p;
	logic landMineExplosion_executed_n;
	logic explosionMineExplosion_executed_p;
	logic explosionMineExplosion_executed_n;
	
	logic [0:15] [0:15] [3:0]  explosionMatrixBitMap_p = '{default:'0}; //don't provide explicit initial values for the array, so it will be initialized with zeroes
	logic [0:15] [0:15] [3:0]  explosionMatrixBitMap_n = '{default:'0};
logic[0:31][0:31][7:0] object_colors = {
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hff,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hde,8'hda,8'hff,8'hff,8'hda,8'hff,8'hda,8'hda,8'hff,8'hda,8'hda,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hff},
	{8'hff,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hda,8'hff,8'hff,8'hf6,8'ha0,8'hff,8'hda,8'hff,8'hff,8'ha0,8'hff,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hda,8'hda,8'hff,8'hda,8'hda,8'hff,8'hda,8'hff},
	{8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hff,8'hff,8'hfa,8'ha0,8'hc4,8'ha0,8'hff,8'hfb,8'hda,8'ha0,8'hfa,8'ha0,8'ha0,8'hfa,8'ha0,8'ha0,8'ha0,8'ha0,8'h80,8'hfb,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hff,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hff,8'hfa,8'ha0,8'ha0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc4,8'hd5,8'hd1,8'hc4,8'hc0,8'hd1,8'hff,8'hda,8'hff,8'hfa,8'hf6,8'hff,8'hff,8'hda,8'hff,8'hff},
	{8'hff,8'hff,8'hda,8'hff,8'hda,8'hda,8'hff,8'h80,8'ha0,8'ha0,8'ha0,8'hc4,8'hcc,8'hcc,8'hcc,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'ha0,8'ha0,8'ha0,8'h80,8'ha0,8'hfa,8'hfa,8'hda,8'hda,8'hff,8'hda,8'hff},
	{8'hff,8'hff,8'hda,8'hff,8'hda,8'hda,8'hcd,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'hcc,8'hcc,8'hcc,8'hf4,8'hc4,8'hc4,8'hcc,8'hcc,8'hc4,8'ha0,8'hc4,8'hc4,8'hc4,8'ha0,8'hfa,8'hda,8'hda,8'hff,8'hda,8'hff},
	{8'hda,8'hff,8'hff,8'h80,8'ha0,8'ha0,8'hc0,8'hc4,8'ha0,8'hc4,8'hd0,8'hd9,8'hd9,8'hd9,8'hd4,8'hcc,8'hcc,8'hcc,8'hcc,8'hec,8'hcc,8'hcc,8'hc4,8'hc4,8'hc4,8'hc4,8'ha0,8'hfe,8'hff,8'hda,8'hff,8'hff},
	{8'hff,8'hff,8'hf6,8'ha0,8'hec,8'hc4,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hd0,8'hd9,8'hd9,8'hd9,8'hd8,8'hd8,8'hd4,8'hf4,8'hf4,8'hc4,8'hc4,8'hcc,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'h80,8'h64,8'hda,8'hff},
	{8'hff,8'hff,8'hf6,8'ha0,8'hcc,8'hec,8'hcc,8'hc4,8'hd4,8'hd4,8'hd0,8'hd4,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd4,8'hf4,8'hcc,8'hcc,8'hcc,8'hcc,8'ha0,8'hc4,8'hc4,8'ha0,8'h60,8'hda,8'hff},
	{8'hda,8'hff,8'hff,8'h80,8'hcc,8'hcc,8'hc4,8'hc4,8'hf4,8'hd4,8'hb0,8'hd9,8'hd9,8'hf9,8'hd4,8'hf9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd4,8'hf4,8'hcc,8'hcc,8'hcc,8'hcc,8'ha0,8'ha0,8'hff,8'hfa,8'hff,8'hff},
	{8'hff,8'hda,8'hda,8'h80,8'hec,8'hcc,8'hcc,8'hcc,8'hd4,8'hd4,8'hd4,8'hf9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd8,8'hd0,8'hcc,8'hc4,8'hcc,8'hc4,8'ha0,8'hfa,8'hff,8'hda,8'hff},
	{8'hff,8'hff,8'hfb,8'h80,8'hc4,8'hcc,8'hcc,8'hcc,8'hd0,8'hd4,8'hd4,8'hd9,8'hd9,8'hd9,8'hd9,8'hfe,8'hff,8'hfe,8'hfe,8'hd9,8'hd9,8'hd8,8'hcc,8'hcc,8'hcc,8'hcc,8'hc4,8'hc4,8'he4,8'h60,8'hda,8'hff},
	{8'ha0,8'ha0,8'hf6,8'he4,8'hc4,8'hcc,8'hcc,8'hcc,8'hcc,8'hd4,8'hd4,8'hd4,8'hd9,8'hd9,8'hfa,8'hff,8'hff,8'hff,8'hff,8'hd9,8'hd9,8'hd4,8'hcc,8'hcc,8'hcc,8'hcc,8'hc4,8'hc4,8'hc4,8'he4,8'hfa,8'hff},
	{8'h80,8'h80,8'hf6,8'hc4,8'hc4,8'hcc,8'hcc,8'hcc,8'hcc,8'hd4,8'hd4,8'hd4,8'hd9,8'hd9,8'hda,8'hff,8'hda,8'hff,8'hfe,8'hd9,8'hd9,8'hd4,8'hcc,8'hec,8'hcc,8'hcc,8'hc4,8'hc4,8'ha0,8'he4,8'hfa,8'hff},
	{8'hff,8'hff,8'hf6,8'hc4,8'hc4,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hd0,8'hd9,8'hd9,8'hfe,8'hfa,8'hff,8'hd9,8'hd9,8'hd9,8'hd9,8'hd4,8'hd4,8'hd4,8'hcc,8'hcc,8'hcc,8'hc4,8'ha0,8'hc4,8'h80,8'hfa,8'hff},
	{8'hda,8'hff,8'hf6,8'he4,8'ha0,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hd0,8'hd4,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd9,8'hd4,8'hd4,8'hd4,8'hc4,8'hc4,8'hcc,8'hc4,8'hc4,8'ha0,8'he4,8'ha0,8'hfa,8'hdf},
	{8'hff,8'hff,8'hda,8'hc4,8'hc4,8'hc4,8'hcc,8'hcc,8'hd4,8'hcc,8'hd4,8'hd4,8'hd4,8'hd4,8'hd8,8'hd9,8'hd9,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd0,8'hcc,8'hcc,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'ha0,8'hff},
	{8'hff,8'hff,8'hf6,8'ha0,8'hc4,8'hc4,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hd0,8'hd4,8'hd4,8'hd0,8'hd0,8'hd0,8'hd4,8'hd4,8'hd4,8'hd4,8'hd0,8'hcc,8'hcc,8'hcc,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'ha0,8'hff},
	{8'hda,8'hff,8'hfa,8'he4,8'hc4,8'hc4,8'hc0,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hd0,8'hd4,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hc4,8'ha0,8'hc4,8'he4,8'ha0,8'hfe},
	{8'hff,8'hff,8'hf6,8'hc4,8'hc4,8'hc4,8'ha0,8'hc4,8'hcc,8'hcc,8'hcc,8'hec,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hc4,8'hc4,8'hc4,8'he4,8'hfa,8'hff},
	{8'hff,8'hff,8'hf6,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'hcc,8'hc4,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hc4,8'hc4,8'hc4,8'ha0,8'h60,8'hda,8'hff},
	{8'hda,8'hff,8'hff,8'h80,8'hc4,8'ha0,8'hc4,8'hc4,8'ha0,8'hc4,8'hc4,8'hcc,8'hcc,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hc4,8'ha0,8'ha0,8'hfa,8'hde,8'hff,8'hff},
	{8'hff,8'hff,8'hda,8'hff,8'ha0,8'ha0,8'ha0,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'hcc,8'hc4,8'hcc,8'hc4,8'hcc,8'hcc,8'he4,8'hfa,8'hda,8'ha0,8'hff,8'hda,8'hff},
	{8'hff,8'hff,8'hda,8'h80,8'hff,8'ha0,8'ha0,8'ha0,8'ha0,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'ha0,8'hc4,8'hc4,8'hc4,8'hc4,8'hcc,8'ha0,8'hc4,8'hc4,8'hc4,8'hfa,8'hfa,8'ha0,8'hff,8'hda,8'hff},
	{8'hda,8'hff,8'hfa,8'hc4,8'hff,8'ha0,8'ha0,8'ha0,8'ha0,8'h80,8'h60,8'h80,8'h80,8'hc4,8'hc4,8'hc4,8'hc4,8'hc4,8'ha0,8'ha0,8'hc4,8'hec,8'hc4,8'he4,8'h60,8'hff,8'h60,8'h60,8'hff,8'hda,8'hff,8'hda},
	{8'hff,8'hff,8'hdf,8'h80,8'ha0,8'hfa,8'hff,8'hff,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hc0,8'hc4,8'hc4,8'hc4,8'hc4,8'ha0,8'ha0,8'hff,8'hff,8'hff,8'hde,8'ha0,8'hfa,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hfa,8'hff,8'hde,8'hda,8'hff,8'hfb,8'hff,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'h80,8'ha0,8'ha0,8'hfa,8'hda,8'hff,8'hff,8'hda,8'hff,8'hda,8'ha0,8'hfa,8'hda,8'hda,8'hff,8'hda,8'hff},
	{8'hda,8'hff,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hda,8'hda,8'hff,8'hda,8'hda,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hff},
	{8'hff,8'hff,8'hda,8'hff,8'hda,8'hda,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hff,8'hda,8'hff,8'hff,8'hff,8'hff,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff}};

 
 
 // pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <= TRANSPARENT_ENCODING ;
	   explosionMatrixBitMap_p = '{default:'0};
		last_direction_p <= 0;
		bombExplosion_executed_p <= 0;
		landMineExplosion_executed_p <= 0;
		explosionMineExplosion_executed_p <= 0;
	end
	else begin
		bombExplosion_executed_p <= bombExplosion_executed_n;
		landMineExplosion_executed_p <= landMineExplosion_executed_n;
		explosionMineExplosion_executed_p <= explosionMineExplosion_executed_n;
		RGBout <= TRANSPARENT_ENCODING ; // default 
		explosionMatrixBitMap_p <= explosionMatrixBitMap_n;
		last_direction_p <= last_direction_n;
		if ((InsideRectangle == 1'b1 )		& 	// only if inside the external bracket 
		   (explosionMatrixBitMap_p[offsetY[8:5] ][offsetX[8:5]] > 4'h0 )) begin // take bits 5,6,7,8,9,10 from address to select  position in the maze    
						RGBout <= object_colors[offsetY[4:0]][offsetX[4:0]] ; 
						if(explosionMatrixBitMap_p[offsetY[8:5] ][offsetX[8:5]] == 4'b0001)
							bombExplosion_executed_p <= 1;
						if(explosionMatrixBitMap_p[offsetY[8:5] ][offsetX[8:5]] == 4'b0010)
							landMineExplosion_executed_p <= 1;
						if(explosionMatrixBitMap_p[offsetY[8:5] ][offsetX[8:5]] == 4'b0100)
							explosionMineExplosion_executed_p <= 1;

		end					
	end 
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
always_comb begin
	last_direction_n = 0;
	explosionMatrixBitMap_n = explosionMatrixBitMap_p;
	bombExplosion_executed_n = bombExplosion_executed_p;
	landMineExplosion_executed_n = landMineExplosion_executed_p;
	explosionMineExplosion_executed_n = explosionMineExplosion_executed_p;
	
	if(explodeBomb && !bombExplosion_executed_p) begin
		last_direction_n = random_dir;
		if(explosionMatrixBitMap_n[bombExplosionIndexY][bombExplosionIndexX] == 0) begin
			case(random_dir ) 
				0: begin //horizontal explosion
							for (int k = 0; k<explosion_length; k++) begin
								if(bombExplosionIndexX+k < 16)
									explosionMatrixBitMap_n[bombExplosionIndexY][bombExplosionIndexX+k] = 4'b0001;
								if(bombExplosionIndexX-k >= 0)	
									explosionMatrixBitMap_n[bombExplosionIndexY][bombExplosionIndexX-k] = 4'b0001; 
							end
					end
				default: begin // vertical explosion
				
						for (int k = 0; k<explosion_length; k++) begin
								if(bombExplosionIndexY+k < 16)
									explosionMatrixBitMap_n[bombExplosionIndexY+k][bombExplosionIndexX] = 4'b0001; 
								if(bombExplosionIndexY-k >= 0)	
									explosionMatrixBitMap_n[bombExplosionIndexY-k][bombExplosionIndexX] = 4'b0001; 
						end
					end
			endcase
		end	
	end
	
	if(mineTriggered && !landMineExplosion_executed_p) begin
		if(explosionMatrixBitMap_n[landMineExplosionIndexY][landMineExplosionIndexY] == 0) begin
			case(random_dir ) 
				0: begin //horizontal explosion
							for (int k = 0; k<explosion_length; k++) begin
								if(landMineExplosionIndexY+k < 16)
									explosionMatrixBitMap_n[landMineExplosionIndexY][landMineExplosionIndexY+k] = 4'b0010; 
								if(landMineExplosionIndexY-k >= 0)	
									explosionMatrixBitMap_n[landMineExplosionIndexY][landMineExplosionIndexY-k] = 4'b0010; 
							end
					end
				default: begin // vertical explosion
				
						for (int k = 0; k<explosion_length; k++) begin
								if(landMineExplosionIndexY+k < 16)
									explosionMatrixBitMap_n[landMineExplosionIndexY+k][explosionMineExplosionIndexX] = 4'b0010; 
								if(landMineExplosionIndexY-k >= 0)	
									explosionMatrixBitMap_n[landMineExplosionIndexY-k][explosionMineExplosionIndexX] = 4'b0010; 
						end
					end
			endcase
		end
	end
	
	
	if(mineExploded && !explosionMineExplosion_executed_p) begin
		case(last_direction_p ) 
			1: begin //horizontal explosion, last direction p = 1 - actual direction ( 1->0, 0->1 )
						for (int k = 0; k<explosion_length; k++) begin
							if(explosionMineExplosionIndexX+k < 16)
								explosionMatrixBitMap_n[explosionMineExplosionIndexY][explosionMineExplosionIndexX+k] = 4'b0100; 
							if(explosionMineExplosionIndexX-k >= 0)	
								explosionMatrixBitMap_n[explosionMineExplosionIndexY][explosionMineExplosionIndexX-k] = 4'b0100; 
						end
				end
			default: begin // vertical explosion
			
					for (int k = 0; k<explosion_length; k++) begin
							if(explosionMineExplosionIndexY+k < 16)
								explosionMatrixBitMap_n[explosionMineExplosionIndexY+k][explosionMineExplosionIndexX] = 4'b0100; 
							if(explosionMineExplosionIndexY-k >= 0)	
								explosionMatrixBitMap_n[explosionMineExplosionIndexY-k][explosionMineExplosionIndexX] = 4'b0100; 
					end
				end
		endcase
	end

		if(OneSecPulse) begin
			for (int i = 0; i <= 15; i++) begin
				for (int j = 0; j <= 15; j++) begin
					if( bombExplosion_executed_p && explosionMatrixBitMap_p[i][j] == 4'b0001) begin
						explosionMatrixBitMap_n[i][j] = 0; //  end explosion
					end 
					if( landMineExplosion_executed_p && explosionMatrixBitMap_p[i][j] == 4'b0010) begin
						explosionMatrixBitMap_n[i][j] = 0; //  end explosion
					end 
					if( explosionMineExplosion_executed_p && explosionMatrixBitMap_p[i][j] == 4'b0100) begin
						explosionMatrixBitMap_n[i][j] = 0; //  end explosion
					end 
				end
			end
			landMineExplosion_executed_n = 0;
			explosionMineExplosion_executed_n = 0;
			bombExplosion_executed_n = 0;
		end	
//		//if ( OneSecPulse ) begin 
//			if(explodeBomb) begin
//				explosionMatrixBitMap_n[bombExplosionIndexY][bombExplosionIndexX] = 4'b0001;
//			end	
//			
//			
//      // Loop through each dimension and initialize to zeroes
//			for (int i = 0; i <= 15; i++) begin
//				for (int j = 0; j <= 15; j++) begin
//						if ( explosionMatrixBitMap_p[i][j] == 4'b0001) begin
//								last_direction_n = random_dir;
//								case(random_dir ) 
//									0: begin //horizontal explosion
//												for (int k = 1; k<explosion_length; k++) begin
//													if(j+k < 16)
//														explosionMatrixBitMap_n[i][j+k] = 4'b0100; // dont put 1 to avoid getting into the if statment
//													if(j-k >= 0)	
//												 		explosionMatrixBitMap_n[i][j-k] = 4'b0100; 
//												end
//										end
//									default: begin // vertical explosion
//									
//											for (int k = 1; k<explosion_length; k++) begin
//													if(i+k < 16)
//														explosionMatrixBitMap_n[i+k][j] = 4'b0100; // dont put 1 to avoid getting into the if statment
//													if(i-k >= 0)	
//														explosionMatrixBitMap_n[i-k][j] = 4'b0100; 
//											end
//										end
//								endcase
//							end // if 2
//						if( explosionMatrixBitMap_p[i][j] > 4'h00) begin
//								explosionMatrixBitMap_n[i][j] = 0; //  end explosion
//						end // if 3
//				end // for 2
//			end // for 1
//		
//		if(mineExploded) begin
//				explosionMatrixBitMap_n[mineExplosionIndexY][mineExplosionIndexX] = 4'b0010;
//		end		
//		
//		for (int i = 0; i <= 15; i++) begin
//				for (int j = 0; j <= 15; j++) begin
//					if ( explosionMatrixBitMap_p[i][j] == 4'b0010) begin
//							case(random_dir ) 
//								0: begin //horizontal explosion
//											for (int k = 1; k<explosion_length; k++) begin
//												if(j+k < 16)
//													explosionMatrixBitMap_n[i][j+k] = 4'b0100; // dont put 1 to avoid getting into the if statment
//												if(j-k >= 0)	
//													explosionMatrixBitMap_n[i][j-k] = 4'b0100; 
//											end
//									end
//								default: begin // vertical explosion
//									
//											for (int k = 1; k<explosion_length; k++) begin
//													if(i+k < 16)
//														explosionMatrixBitMap_n[i+k][j] = 4'b0100; // dont put 1 to avoid getting into the if statment
//													if(i-k >= 0)	
//														explosionMatrixBitMap_n[i-k][j] = 4'b0100; 
//											end
//									end
//							endcase
//					end // if 2
//					if( explosionMatrixBitMap_p[i][j] > 4'h00) begin
//							explosionMatrixBitMap_n[i][j] = 0; //  end explosion
//					end // if 3
//				end
//			end
//			
//			if(mineTriggered) begin
//				explosionMatrixBitMap_n[mineExplosionIndexY][mineExplosionIndexX] = 4'b0011;
//			end
//			
//			for (int i = 0; i <= 15; i++) begin
//				for (int j = 0; j <= 15; j++) begin
//					if ( explosionMatrixBitMap_p[i][j] == 4'b0011) begin
//										case(last_direction_p ) 
//											0: begin //horizontal explosion
//														for (int k = 1; k<explosion_length; k++) begin
//															if(j+k < 16)
//																explosionMatrixBitMap_n[i][j+k] = 4'b0100; // dont put 3 to avoid getting into the if statment
//															if(j-k >= 0)	
//																explosionMatrixBitMap_n[i][j-k] = 4'b0100; 
//														end
//												end
//											default: begin // vertical explosion
//											
//													for (int k = 1; k<explosion_length; k++) begin
//															if(i+k < 16)
//																explosionMatrixBitMap_n[i+k][j] = 4'b0100; // dont put 3 to avoid getting into the if statment
//															if(i-k >= 0)	
//																explosionMatrixBitMap_n[i-k][j] = 4'b0100; 
//													end
//												end
//										endcase
//									end
//						if( explosionMatrixBitMap_p[i][j] > 4'b0000) begin
//								explosionMatrixBitMap_n[i][j] = 0; //  end explosion
//						end // if 3
//				end // for 2
//			end
			
end // start comb
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule

