// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen Apr  2023  
// (c) Technion IIT, Department of Electrical Engineering 2023 



module	wallMatrixBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input logic wall_explode,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic OneSecPulse,
					
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout,  //rgb value from the bitmap 
					output logic increase_score
 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */

// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 16*16 and use only the top left 16*15 squares 
// this is the bitmap  of the maze , if there is a specific value  the  whole 32*32 rectange will be drawn on the screen
// there are  16 options of differents kinds of 32*32 squares 
// all numbers here are hard coded to simplify the  understanding 
// wall_4 -> blue (unbreakable)
// wall_3 -> grey
// wall_2 -> brown
// wall_1 -> yellow
logic explosion_executed_p = 0;
logic explosion_executed_n = 0;
const logic [0:31][0:31][7:0] wall_4 = {
	{8'h04,8'h2d,8'h04,8'h04,8'h0d,8'h04,8'h04,8'h0d,8'h2d,8'h04,8'h0d,8'h0d,8'h04,8'h32,8'h72,8'h9b,8'h04,8'h72,8'h72,8'h72,8'h72,8'h9b,8'h04,8'h0d,8'h72,8'h72,8'h76,8'h05,8'h04,8'h04,8'h04,8'h0d},
	{8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h04,8'h0d,8'h72,8'h9b,8'h0d,8'h72,8'h72,8'h72,8'h72,8'h32,8'h04,8'h0d,8'h72,8'h72,8'h9b,8'h05,8'h9b,8'h32,8'h9b,8'h9b},
	{8'h72,8'h9b,8'h0d,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h32,8'h2d,8'h72,8'h72,8'h9b,8'h04,8'h0d,8'h72,8'h72,8'h72,8'h9b,8'h04,8'h2d,8'h72,8'h72,8'h9b,8'h05,8'h32,8'h32,8'h72,8'h32},
	{8'h2d,8'h9f,8'h05,8'h0d,8'h2d,8'h2d,8'h2d,8'h0d,8'h2d,8'h0d,8'h2d,8'h2d,8'h04,8'h2d,8'h2d,8'h2e,8'h0d,8'h72,8'h72,8'h72,8'h72,8'h72,8'h04,8'h72,8'h72,8'h72,8'h72,8'h05,8'h0d,8'h2d,8'h0d,8'h2d},
	{8'h0e,8'h9b,8'h9b,8'hbb,8'h04,8'h2d,8'h04,8'h04,8'h04,8'h04,8'h04,8'h04,8'h04,8'h04,8'h32,8'h9b,8'h05,8'h2e,8'h72,8'h0d,8'h0d,8'h9f,8'h04,8'h0e,8'h72,8'h72,8'hbf,8'h05,8'h9b,8'h9b,8'h9b,8'hbf},
	{8'h0d,8'h32,8'h72,8'h76,8'h9b,8'h72,8'h72,8'h72,8'h04,8'h72,8'h32,8'h72,8'h04,8'h04,8'h04,8'h2e,8'h0d,8'h05,8'h05,8'h05,8'h05,8'h2d,8'h04,8'h05,8'h0e,8'h05,8'h05,8'h04,8'h72,8'h32,8'h72,8'h9b},
	{8'h2e,8'h72,8'h72,8'h32,8'h9b,8'h32,8'h72,8'h72,8'h72,8'h32,8'h72,8'h72,8'h72,8'h04,8'h9b,8'h9b,8'h9b,8'h9b,8'h2e,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h04,8'h05,8'h72,8'h72,8'h9b},
	{8'h04,8'h0d,8'h72,8'h32,8'hbb,8'h72,8'h72,8'h72,8'h32,8'h72,8'h32,8'h72,8'h72,8'h04,8'h0d,8'h72,8'h72,8'h32,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h32,8'h72,8'h72,8'h05,8'h72,8'h72,8'h72,8'h72},
	{8'h05,8'h0d,8'h32,8'h32,8'hbb,8'h72,8'h72,8'h9b,8'h9b,8'h72,8'h9b,8'h32,8'h72,8'h05,8'h2d,8'h72,8'h72,8'h32,8'h32,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h9b,8'h05,8'h05,8'h04,8'h72,8'h9b},
	{8'h04,8'h04,8'h04,8'h05,8'h04,8'h72,8'h72,8'h04,8'h04,8'h72,8'h72,8'h72,8'h04,8'h04,8'h0d,8'h72,8'h72,8'h0d,8'h72,8'h72,8'h72,8'h9b,8'h32,8'h72,8'h72,8'h72,8'h72,8'h04,8'h0d,8'h05,8'h32,8'h9b},
	{8'h2e,8'h72,8'h72,8'hbb,8'h32,8'h9b,8'h72,8'h9b,8'h2e,8'h72,8'h72,8'h72,8'h72,8'h9b,8'h2d,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h32,8'h0e,8'h0d,8'h0d,8'h72,8'h9b},
	{8'h04,8'h0d,8'h2d,8'hbb,8'h2d,8'h72,8'h72,8'h9b,8'h04,8'h2d,8'h0d,8'h0d,8'h2d,8'h9b,8'h2d,8'h2d,8'h0d,8'h2d,8'h2d,8'h0d,8'h2d,8'h2d,8'h32,8'h0e,8'h2d,8'h2d,8'h2d,8'h05,8'h0d,8'h0d,8'h05,8'h04},
	{8'h9b,8'h9b,8'h9b,8'hbb,8'h2e,8'h72,8'h72,8'h9b,8'h0d,8'h9b,8'h9b,8'h9b,8'hbf,8'h9b,8'h9b,8'h9b,8'h0e,8'h9b,8'hbb,8'h9b,8'h32,8'h9b,8'hbb,8'h9b,8'h9b,8'h0e,8'h9b,8'hbf,8'h32,8'h9b,8'h9b,8'h9b},
	{8'h76,8'h72,8'h72,8'hbb,8'h2e,8'h2e,8'h2e,8'h9b,8'h05,8'h32,8'h72,8'h9b,8'h2d,8'h32,8'h72,8'h9b,8'h05,8'h72,8'h32,8'h72,8'h72,8'h72,8'h32,8'h72,8'h9b,8'h04,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h72,8'h72,8'h32,8'h72,8'h05,8'h05,8'h05,8'h05,8'h04,8'h72,8'h72,8'h9b,8'h2d,8'h72,8'h72,8'h9b,8'h04,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h9b,8'h2d,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h0e,8'h04,8'h0d,8'hbb,8'h72,8'h72,8'h32,8'h32,8'h2d,8'h72,8'h72,8'h32,8'h0d,8'h05,8'h72,8'h9b,8'h04,8'h72,8'h72,8'h2e,8'h72,8'h72,8'h72,8'h72,8'h9b,8'h04,8'h0d,8'h2d,8'h2d,8'h0d,8'h0d,8'h0d},
	{8'h32,8'h9b,8'hbb,8'h04,8'h04,8'h04,8'h04,8'h04,8'h04,8'h72,8'h32,8'h9b,8'h04,8'h2e,8'h72,8'h9b,8'h04,8'h0d,8'h0d,8'h72,8'h2d,8'h72,8'h72,8'h0d,8'h9b,8'h9b,8'h9b,8'h72,8'h72,8'h9b,8'h9b,8'h9b},
	{8'hbb,8'h72,8'hbb,8'hbb,8'h72,8'h72,8'h72,8'h05,8'h05,8'h2e,8'h0d,8'h0e,8'h05,8'h0d,8'h0d,8'h2d,8'h04,8'h04,8'h04,8'h04,8'h04,8'h04,8'h04,8'h04,8'h04,8'h0d,8'h72,8'h32,8'h32,8'h72,8'h72,8'h32},
	{8'h72,8'h72,8'h72,8'h32,8'h72,8'h2e,8'h72,8'h05,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'hbb,8'h9b,8'h32,8'h9b,8'h2e,8'h0d,8'h05,8'h05,8'h72,8'h05,8'h05,8'h05,8'h04,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72},
	{8'h0d,8'h72,8'hbb,8'h9b,8'h32,8'h9b,8'h32,8'h0d,8'h04,8'h32,8'h72,8'h72,8'h72,8'h72,8'h72,8'h9b,8'h9b,8'h32,8'h32,8'h32,8'h72,8'h2e,8'h72,8'h72,8'h0e,8'h05,8'h2d,8'h2d,8'h0d,8'h0d,8'h72,8'h72},
	{8'h2d,8'hbb,8'hbb,8'h2d,8'h05,8'hbb,8'h72,8'h9b,8'h04,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h9b,8'h9b,8'h9b,8'h32,8'h2d,8'hbb,8'h9b,8'h2e,8'hbb,8'h9b,8'hbb,8'h72,8'hbb,8'hbb,8'h2d,8'hbb,8'hbb},
	{8'h9b,8'h32,8'h72,8'h32,8'h0d,8'h32,8'h32,8'h9b,8'h0d,8'h05,8'h72,8'h72,8'h72,8'h72,8'h72,8'h9b,8'h0e,8'h32,8'h32,8'h9b,8'h0d,8'h72,8'h9b,8'h32,8'h72,8'h32,8'hbb,8'h2e,8'h32,8'h77,8'h32,8'h32},
	{8'h0d,8'h72,8'h0d,8'h72,8'h05,8'h32,8'h72,8'h9b,8'h0d,8'h0d,8'h04,8'h05,8'h72,8'h72,8'h72,8'h9b,8'h04,8'h72,8'h72,8'h9b,8'h05,8'h72,8'h72,8'h72,8'h72,8'h72,8'h9b,8'h04,8'h72,8'h72,8'h0d,8'h72},
	{8'h04,8'h04,8'h05,8'h04,8'h04,8'h04,8'h04,8'h04,8'h32,8'h0d,8'h04,8'h04,8'h72,8'h72,8'h72,8'h9b,8'h04,8'h2e,8'h72,8'hbb,8'h0e,8'h32,8'h72,8'h72,8'h72,8'h72,8'h9b,8'h04,8'h04,8'h04,8'h04,8'h04},
	{8'h0d,8'h04,8'h72,8'h0d,8'h05,8'h04,8'h0d,8'h04,8'h72,8'h0d,8'h2d,8'h72,8'h72,8'h72,8'h72,8'h72,8'h2d,8'h72,8'h72,8'h9b,8'h0d,8'h72,8'h72,8'h72,8'h72,8'h9b,8'h32,8'h9b,8'h04,8'h04,8'h2d,8'h04},
	{8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h04,8'h32,8'h0d,8'h0d,8'h05,8'h04,8'h0e,8'h05,8'h04,8'h0d,8'h72,8'h72,8'hbb,8'h2d,8'h72,8'h72,8'h72,8'h72,8'h72,8'h9b,8'h9b,8'h32,8'h72,8'h72,8'h32},
	{8'h72,8'h72,8'h32,8'h72,8'h72,8'h72,8'h72,8'h04,8'h0e,8'h2e,8'h05,8'h05,8'hbf,8'h9b,8'h32,8'h9b,8'h04,8'h72,8'h72,8'h9b,8'h04,8'h72,8'h72,8'h72,8'h72,8'h32,8'h72,8'h9b,8'h72,8'h72,8'h2e,8'h72},
	{8'h9b,8'h32,8'h32,8'h32,8'h32,8'h32,8'h72,8'h05,8'h9f,8'h72,8'h2e,8'h72,8'h2d,8'h32,8'h9b,8'h9b,8'h0d,8'h72,8'h32,8'h9b,8'h0d,8'h72,8'h72,8'h0d,8'h72,8'h72,8'h9f,8'h9b,8'h77,8'h32,8'h72,8'h32},
	{8'h05,8'h32,8'h32,8'h72,8'h72,8'h32,8'h32,8'h72,8'h05,8'h05,8'h05,8'h05,8'h04,8'h32,8'h72,8'h9b,8'h04,8'h05,8'h04,8'h04,8'h04,8'h05,8'h05,8'h04,8'h05,8'h04,8'h05,8'h05,8'h32,8'h32,8'h05,8'h72},
	{8'h9b,8'h32,8'h05,8'h32,8'h9b,8'h72,8'h9b,8'h9b,8'h32,8'h9b,8'h32,8'h32,8'h2d,8'h0d,8'h72,8'h9b,8'h0d,8'h32,8'h9b,8'h9b,8'h32,8'h9b,8'h05,8'h32,8'h9b,8'h32,8'h72,8'h05,8'h32,8'h9b,8'h9b,8'h9b},
	{8'h32,8'h32,8'h05,8'h0d,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h32,8'h2d,8'h0d,8'h72,8'h9b,8'h05,8'h2e,8'h72,8'h72,8'h72,8'h9b,8'h04,8'h2e,8'h72,8'h72,8'h9b,8'h04,8'h32,8'h72,8'h72,8'h72},
	{8'h72,8'h9b,8'h05,8'h2d,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h9b,8'h04,8'h72,8'h72,8'h9b,8'h0d,8'h72,8'h72,8'h72,8'h72,8'h72,8'h05,8'h0e,8'h72,8'h72,8'h9b,8'h05,8'h0d,8'h72,8'h72,8'h72}
	};


const logic [0:31][0:31][7:0] wall_3 = {
	{8'hb6,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'hb6,8'hb6,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h96,8'h95,8'h96,8'h91,8'hb6,8'hb2,8'h91,8'h95,8'h92,8'hb6,8'hb6,8'hb6,8'h91},
	{8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h24,8'h00,8'h25,8'h92,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h96,8'h2d,8'h24,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'h92,8'hff},
	{8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h71,8'h92,8'h91,8'h24,8'h92,8'h92,8'h92,8'h92,8'h96,8'h6d,8'h6d,8'h92,8'h92,8'h92,8'h92,8'h6d,8'h6d,8'h6d,8'h71,8'h91,8'h24,8'h96,8'h96,8'h71,8'h71,8'h6d,8'hff},
	{8'hb6,8'hb6,8'hb6,8'hb6,8'h92,8'h92,8'h92,8'h91,8'h24,8'h96,8'h96,8'h91,8'h91,8'h91,8'h6d,8'h6d,8'h91,8'h91,8'h91,8'h91,8'h6d,8'h71,8'h71,8'h6d,8'h6d,8'h24,8'h71,8'h71,8'h71,8'h71,8'h71,8'hff},
	{8'hb6,8'hb6,8'h91,8'h91,8'h91,8'h92,8'h92,8'h6d,8'h24,8'h92,8'h6d,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h91,8'h6d,8'h6d,8'h6d,8'h71,8'h71,8'h6d,8'h6d,8'h24,8'h71,8'h6d,8'h71,8'h71,8'h71,8'hff},
	{8'hb6,8'hb6,8'h91,8'h91,8'h91,8'h92,8'h6d,8'h6d,8'h24,8'h96,8'h71,8'h71,8'h71,8'h91,8'h6d,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h8d,8'h71,8'h71,8'h6d,8'h6d,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hff},
	{8'hb6,8'hb6,8'h92,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h96,8'h6d,8'h71,8'h6d,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h91,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h71,8'h6d,8'h6d,8'h71,8'h8d,8'hff},
	{8'hb6,8'hb6,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h6d,8'h6d,8'h71,8'h6d,8'h65,8'hff},
	{8'hb6,8'hb6,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h25,8'h65,8'h6d,8'h6d,8'h65,8'hff},
	{8'hb6,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h24,8'hff},
	{8'hb6,8'h24,8'h92,8'hb6,8'h96,8'h96,8'h96,8'h96,8'h96,8'h96,8'h24,8'h91,8'h91,8'h91,8'h71,8'h71,8'h91,8'h71,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'hb6,8'hb6,8'h92,8'h00,8'h24,8'hff},
	{8'hb6,8'hb6,8'h71,8'h6d,8'h71,8'hb6,8'h96,8'h71,8'h6d,8'h6d,8'h6d,8'h91,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h25,8'h24,8'h96,8'h96,8'h6d,8'h92,8'h96,8'h92,8'h6d,8'h6d,8'h6d,8'h71,8'h91,8'hff},
	{8'hb6,8'hb6,8'h71,8'h6d,8'h6d,8'h96,8'h96,8'h6d,8'h6d,8'h6d,8'h6d,8'h71,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h25,8'h24,8'h96,8'h96,8'h6d,8'h92,8'hb6,8'hb6,8'h6d,8'h6d,8'h71,8'h6d,8'h91,8'hff},
	{8'hb6,8'hb6,8'h91,8'h71,8'h6d,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h25,8'h24,8'h96,8'h6d,8'h91,8'h6d,8'h6d,8'h71,8'h91,8'h91,8'h91,8'h6d,8'h6d,8'hff},
	{8'hb6,8'hb6,8'h6d,8'h6d,8'h65,8'h65,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h25,8'h25,8'h25,8'h25,8'h25,8'h24,8'h6d,8'h6d,8'h71,8'h6d,8'h65,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hff},
	{8'hb6,8'hb6,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h2d,8'h25,8'h2d,8'h25,8'h25,8'h25,8'h25,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hff},
	{8'hb6,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'hff},
	{8'hb6,8'hb6,8'h96,8'hb6,8'h24,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h04,8'h24,8'h92,8'h96,8'h96,8'h92,8'h92,8'h92,8'h96,8'hb6,8'hff},
	{8'hb6,8'hb6,8'h91,8'h91,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'h92,8'h91,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h91,8'h91,8'h92,8'h92,8'h6d,8'h24,8'h92,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h91,8'h91,8'h91,8'hff},
	{8'hb6,8'hb6,8'h91,8'h6d,8'h24,8'hb6,8'hb6,8'h92,8'h92,8'h92,8'h92,8'h91,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h92,8'h92,8'h6d,8'h8d,8'h24,8'h96,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h91,8'h91,8'h91,8'hff},
	{8'hb6,8'hb6,8'h6d,8'h6d,8'h24,8'h92,8'h92,8'h92,8'h6d,8'h6d,8'h92,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h8d,8'h6d,8'h24,8'h6d,8'h6d,8'h6d,8'h25,8'h25,8'h65,8'h65,8'h65,8'h25,8'hff},
	{8'hb6,8'hb6,8'h6d,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h65,8'h25,8'h65,8'h25,8'h25,8'h65,8'h65,8'h65,8'h25,8'hff},
	{8'hb6,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h71,8'h96,8'h96,8'h96,8'h96,8'h92,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'hff},
	{8'hb6,8'h91,8'h96,8'h96,8'h96,8'h96,8'h96,8'h96,8'h96,8'h96,8'h92,8'h71,8'h71,8'h91,8'h96,8'h96,8'h96,8'h96,8'h96,8'h96,8'h71,8'h91,8'h6d,8'h6d,8'h6d,8'h91,8'h6d,8'h6d,8'h6d,8'h25,8'h6d,8'hff},
	{8'hb6,8'hb6,8'h96,8'h96,8'h96,8'h96,8'h96,8'h96,8'h96,8'h92,8'h71,8'h71,8'h6d,8'h71,8'hb6,8'h96,8'hb6,8'h96,8'h96,8'hb6,8'h6d,8'h71,8'h6d,8'h91,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hff},
	{8'hb6,8'hb6,8'h96,8'h91,8'h91,8'h71,8'h96,8'h96,8'h71,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'hb6,8'h96,8'h71,8'h96,8'h92,8'h6d,8'h6d,8'h6d,8'h25,8'h71,8'h92,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hff},
	{8'hb6,8'hb6,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'hb6,8'h92,8'h6d,8'h6d,8'h6d,8'h6d,8'h91,8'h2d,8'h6d,8'h71,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h25,8'h25,8'hff},
	{8'hb6,8'hb6,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'hb6,8'h92,8'h6d,8'h6d,8'h71,8'h6d,8'h91,8'h65,8'h6d,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h25,8'hff},
	{8'hb6,8'hb6,8'h71,8'h71,8'h65,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h65,8'h6d,8'h6d,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'hff},
	{8'hb6,8'h00,8'h6d,8'h6d,8'h65,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h65,8'h24,8'h24,8'h25,8'h65,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h6d,8'h65,8'h25,8'h25,8'h25,8'h24,8'h24,8'hff},
	{8'hb6,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h65,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h25,8'h25,8'h25,8'h25,8'h24,8'h24,8'h24,8'hff},
	{8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff}
	};
const logic [0:31][0:31][7:0] wall_2 = {
	{8'h24,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h24,8'h20,8'h20,8'h24,8'h64,8'h64,8'h64,8'h64,8'h24,8'h64,8'h64,8'h24,8'h20,8'h64,8'h64,8'h20,8'h24,8'h20,8'h24,8'h24,8'h64,8'h6d,8'h6d,8'h24,8'h64},
	{8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'hd6,8'h91,8'hb1,8'hfa,8'hd5,8'hd5,8'hd6,8'hd6,8'h20,8'hd6,8'h91,8'h91,8'h91,8'hb5,8'h64,8'h20,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb5,8'h91,8'h00,8'h64,8'h6d},
	{8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h20,8'hb1,8'hb1,8'h91,8'hb1,8'hb1,8'h64,8'h20,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h20,8'h64,8'h64},
	{8'h20,8'h24,8'h20,8'h24,8'h20,8'h20,8'h20,8'h24,8'h24,8'h20,8'h20,8'h24,8'h20,8'h00,8'h00,8'h24,8'h64,8'h24,8'h64,8'h24,8'h00,8'h24,8'h20,8'h24,8'h64,8'h6c,8'h20,8'h20,8'h00,8'h20,8'h20,8'h20},
	{8'h20,8'h20,8'hd5,8'hd5,8'hb5,8'hd5,8'hb5,8'hb1,8'h91,8'h20,8'hda,8'hb1,8'h91,8'hd5,8'hd5,8'h20,8'hb1,8'h6c,8'h91,8'h91,8'hb1,8'hb5,8'h6c,8'h64,8'h8d,8'h20,8'hb5,8'hd5,8'hb5,8'hb1,8'hb1,8'hb1},
	{8'h24,8'h20,8'h8c,8'hb1,8'hb1,8'hb1,8'h91,8'hb1,8'h91,8'h64,8'hb1,8'h8d,8'h91,8'h91,8'hb1,8'h64,8'h8d,8'h8c,8'hb1,8'hb1,8'h6c,8'h6c,8'h6c,8'h6c,8'h8d,8'h00,8'h8d,8'h8d,8'h8d,8'h8d,8'h8c,8'h8d},
	{8'h64,8'h24,8'h8c,8'h91,8'h91,8'h91,8'h91,8'h91,8'h8d,8'h00,8'h8d,8'h91,8'h91,8'h91,8'h91,8'h20,8'h64,8'h6d,8'h64,8'h91,8'h6c,8'h6c,8'h6c,8'h6c,8'h64,8'h20,8'h8d,8'h6c,8'h8c,8'h8c,8'h6c,8'h6c},
	{8'h6d,8'h20,8'hb1,8'h8d,8'h91,8'h6c,8'h24,8'h6c,8'h24,8'h00,8'h91,8'h91,8'h91,8'h91,8'hb1,8'h20,8'h64,8'h64,8'h20,8'h24,8'h6c,8'h6c,8'h6c,8'h6c,8'h64,8'h20,8'h8c,8'h6c,8'h6c,8'h6c,8'h6c,8'h6c},
	{8'h20,8'h20,8'h20,8'h64,8'h64,8'h00,8'h20,8'h20,8'h24,8'h20,8'h20,8'h24,8'h64,8'h64,8'h6c,8'h24,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h6c,8'h8d,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20},
	{8'h64,8'h64,8'h64,8'h64,8'h64,8'h24,8'h8c,8'h8c,8'h6c,8'h6c,8'h8c,8'h8c,8'h6c,8'h64,8'h8d,8'h91,8'h91,8'h91,8'h91,8'h91,8'hd6,8'h8c,8'h91,8'h91,8'h91,8'h91,8'h8d,8'h8c,8'h8d,8'h20,8'h64,8'h64},
	{8'h64,8'h64,8'h64,8'h24,8'h20,8'h20,8'h64,8'h8c,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h20,8'h8d,8'h8d,8'h91,8'hb1,8'h91,8'h91,8'h91,8'h91,8'h91,8'h8d,8'h8d,8'h8d,8'h8d,8'h91,8'h91,8'h00,8'h24,8'h64},
	{8'h64,8'h64,8'h24,8'h24,8'h20,8'h20,8'h24,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h24,8'h24,8'h00,8'h20,8'h24,8'h24,8'h20,8'h6c,8'h6c,8'h8d,8'h91,8'h91,8'h8d,8'h91,8'h91,8'h00,8'h20,8'h20},
	{8'h20,8'h20,8'h91,8'hb1,8'hb1,8'h8d,8'h20,8'h20,8'h20,8'h8d,8'h8d,8'h00,8'hfa,8'h8d,8'h91,8'h24,8'hb1,8'hd5,8'hd5,8'hb5,8'hb1,8'h00,8'h20,8'h00,8'h20,8'hb1,8'hb1,8'h24,8'h8d,8'h6c,8'h91,8'h91},
	{8'h91,8'h64,8'hd5,8'hb1,8'h91,8'h8c,8'h91,8'h00,8'h91,8'h91,8'h91,8'h24,8'h8d,8'h8d,8'h91,8'h91,8'h91,8'h8d,8'h8d,8'h91,8'hb1,8'hd5,8'hb5,8'h20,8'h6c,8'h6c,8'h64,8'h6d,8'h6c,8'h8c,8'h6c,8'h8c},
	{8'h64,8'h24,8'hb1,8'h91,8'h8d,8'h91,8'h8d,8'h24,8'hb1,8'h91,8'h91,8'h20,8'h20,8'h20,8'h6d,8'h91,8'h8d,8'h8d,8'h8d,8'h8d,8'h91,8'h91,8'h8d,8'h20,8'h6d,8'h64,8'h64,8'h64,8'h6c,8'h8d,8'h6c,8'h6c},
	{8'h24,8'h64,8'hb1,8'h8d,8'h91,8'h91,8'hb5,8'h64,8'h8d,8'h91,8'hb1,8'h24,8'hb1,8'hb1,8'hb1,8'h64,8'h91,8'h8d,8'h8d,8'h8d,8'hb1,8'h64,8'h64,8'h20,8'h6c,8'h24,8'h64,8'h20,8'h24,8'h6c,8'h64,8'h6c},
	{8'h20,8'h20,8'h24,8'h8d,8'h6d,8'h6d,8'h24,8'h24,8'h20,8'h24,8'h64,8'h20,8'h24,8'h64,8'h6d,8'h00,8'h64,8'h20,8'h24,8'h24,8'h20,8'h24,8'hb1,8'h91,8'h6d,8'h64,8'h64,8'h64,8'h24,8'h24,8'h20,8'h20},
	{8'h8d,8'h91,8'hb1,8'hd5,8'hd5,8'h20,8'hb5,8'h8c,8'h8c,8'h64,8'h91,8'hb1,8'h6c,8'h20,8'h20,8'h6d,8'h64,8'h6d,8'h64,8'h20,8'hb1,8'h8c,8'h8c,8'h8c,8'h64,8'h64,8'h64,8'h20,8'h8d,8'h91,8'h91,8'hb1},
	{8'hb1,8'hb1,8'h8d,8'hb1,8'h91,8'h20,8'hd5,8'h8c,8'h8c,8'h64,8'h8c,8'h6c,8'h6c,8'h24,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h6d,8'h6c,8'h6c,8'h6c,8'h8c,8'h64,8'h64,8'h64,8'h24,8'h8d,8'hb1,8'h91,8'h91},
	{8'h91,8'h91,8'hb1,8'h91,8'hb1,8'h24,8'h8d,8'h8c,8'h6c,8'h20,8'h64,8'h24,8'h64,8'h24,8'h24,8'h24,8'h20,8'h24,8'h24,8'h24,8'h64,8'h64,8'h6c,8'h6c,8'h64,8'h00,8'h20,8'h20,8'h20,8'h64,8'h91,8'h91},
	{8'h91,8'h20,8'h6d,8'h8d,8'h8d,8'h64,8'h64,8'h8c,8'h6c,8'hb1,8'h91,8'h91,8'h91,8'hb1,8'hb1,8'h6c,8'hd6,8'h91,8'h64,8'hb1,8'h91,8'hb1,8'hb1,8'h91,8'hb1,8'hb1,8'h24,8'h91,8'h91,8'h91,8'h91,8'h91},
	{8'h6c,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h6c,8'hb1,8'h91,8'h91,8'h91,8'h91,8'hb1,8'h24,8'h24,8'hb1,8'h64,8'h6c,8'h91,8'h91,8'h8d,8'h91,8'h8d,8'hb1,8'h24,8'h91,8'h8d,8'h8d,8'h91,8'h91},
	{8'h24,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h8c,8'hb5,8'h91,8'h91,8'h64,8'h91,8'h91,8'h64,8'h20,8'h24,8'h24,8'h20,8'h24,8'h24,8'h64,8'h64,8'h91,8'h00,8'h00,8'h91,8'h8d,8'h8d,8'hb1,8'h91},
	{8'h20,8'h65,8'h64,8'h64,8'h24,8'h64,8'h24,8'h20,8'h24,8'hb5,8'hb1,8'h91,8'h91,8'h64,8'h64,8'h20,8'hb5,8'hd5,8'hd5,8'h20,8'h24,8'h24,8'h24,8'h64,8'h24,8'h00,8'h20,8'h20,8'h24,8'h24,8'h20,8'h20},
	{8'hd5,8'h91,8'h91,8'h00,8'h00,8'h20,8'h24,8'hb5,8'hb1,8'h00,8'h20,8'h24,8'h00,8'h00,8'h24,8'h91,8'h91,8'hb1,8'hb5,8'h8d,8'h20,8'h20,8'h20,8'h20,8'h6c,8'h6c,8'h6c,8'h91,8'h91,8'h20,8'hd5,8'hb5},
	{8'h91,8'h91,8'hb1,8'h91,8'h91,8'h8d,8'h64,8'h8c,8'h8d,8'h6c,8'h6c,8'h6c,8'h6c,8'h6c,8'h8c,8'h24,8'h91,8'h91,8'h64,8'hb1,8'h91,8'h91,8'h20,8'h64,8'h91,8'h8d,8'h8d,8'h91,8'h91,8'h20,8'h91,8'h91},
	{8'h91,8'hb1,8'hb1,8'h91,8'h8d,8'h6d,8'h20,8'h91,8'h64,8'h8d,8'h8c,8'h8d,8'h8d,8'h20,8'h8d,8'h24,8'hb5,8'h91,8'hb1,8'h24,8'h8d,8'hb1,8'h20,8'h24,8'h64,8'h24,8'h8d,8'h64,8'h64,8'h24,8'hb1,8'hb1},
	{8'h64,8'h64,8'h64,8'h64,8'h64,8'h00,8'h6c,8'h64,8'h24,8'h20,8'h20,8'h20,8'h64,8'h64,8'h6d,8'h24,8'h20,8'h64,8'h00,8'hd5,8'h24,8'h20,8'h20,8'h20,8'h24,8'h00,8'h20,8'h24,8'h24,8'h24,8'h6d,8'h64},
	{8'h20,8'h91,8'hb5,8'hb5,8'h8c,8'h6c,8'h8c,8'h6c,8'h6c,8'h20,8'hb1,8'h91,8'hb1,8'h24,8'h64,8'hb5,8'hd5,8'hfa,8'h20,8'h91,8'h6c,8'h8d,8'h8c,8'hb1,8'hb1,8'h64,8'hb1,8'h91,8'h91,8'hb1,8'h8d,8'h24},
	{8'h24,8'hb5,8'h6c,8'h8d,8'h6c,8'h8d,8'h64,8'h6c,8'h8d,8'h00,8'h91,8'h91,8'h24,8'h24,8'h91,8'h91,8'hb1,8'h91,8'h20,8'hb1,8'h8c,8'h8c,8'h8c,8'h8d,8'h64,8'h6c,8'h91,8'h8d,8'h91,8'h8d,8'h8d,8'h91},
	{8'h64,8'h91,8'h8c,8'h8d,8'h6c,8'h6c,8'h6c,8'h6c,8'h6c,8'h20,8'h6c,8'h24,8'hb5,8'h91,8'h91,8'h91,8'h91,8'h91,8'h24,8'hb1,8'h6c,8'h8c,8'h8c,8'h6c,8'h24,8'h24,8'h91,8'h91,8'h91,8'h91,8'hb1,8'h91},
	{8'h8d,8'h6c,8'h64,8'h6c,8'h6c,8'h6c,8'h6c,8'h6c,8'h8c,8'h24,8'hb5,8'h91,8'h91,8'hb1,8'h91,8'h91,8'h91,8'hb1,8'h6c,8'h64,8'h6c,8'h6c,8'h64,8'h8d,8'h64,8'h64,8'h91,8'h91,8'h91,8'h8d,8'h8d,8'h91}
	};
const logic [0:31][0:31][7:0] wall_1 = {
	{8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hf9,8'hf0,8'hf4,8'hf8,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf0,8'hf8,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe},
	{8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hf9,8'hf4,8'hf8,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hf9,8'hfe,8'hfd,8'hf8,8'hfc,8'hfd,8'hf0,8'hf9,8'hf9,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe},
	{8'hf9,8'hfd,8'hfe,8'hfe,8'hf9,8'hf9,8'hf0,8'hf9,8'hf9,8'hfd,8'hfd,8'hf9,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hf8,8'hfd,8'hf8,8'hf4,8'hf0,8'hf9,8'hfd,8'hf9,8'hf9,8'hfd},
	{8'hfd,8'hf9,8'hf0,8'hf0,8'hf9,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hf9,8'hfd,8'hfd,8'hf9,8'hfd,8'hf9,8'hfd,8'hf9,8'hfd},
	{8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hf9,8'hfd,8'hfd,8'hfe,8'hf9,8'hfd,8'hfd},
	{8'hfe,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfe,8'hfd,8'hfe,8'hfe},
	{8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe},
	{8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe},
	{8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe},
	{8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hf8,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe},
	{8'hfe,8'hfd,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hfd,8'hfd,8'hf4,8'hf4,8'hf4,8'hf4,8'hfd,8'hf4,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe},
	{8'hf4,8'hf8,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf8,8'hf9,8'hf4,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd},
	{8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfd,8'hfd,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hfd,8'hfd,8'hfd,8'hfd,8'hf0,8'hf9,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hf9,8'hf0,8'hf9},
	{8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf0,8'hf0,8'hf0,8'hf0,8'hf9,8'hf9,8'hf9,8'hfd},
	{8'hfd,8'hfd,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe},
	{8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hf9,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hf9,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe},
	{8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfd,8'hfe},
	{8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe},
	{8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe},
	{8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hf9,8'hf0,8'hf0,8'hf0,8'hf0,8'hf4,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe},
	{8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hf0,8'hf8,8'hfd,8'hfd,8'hfd,8'hfe,8'hf9,8'hf0,8'hf4,8'hf9,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfe},
	{8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hf4,8'hfd,8'hf9,8'hfd,8'hfd,8'hfd,8'hfe,8'hfd,8'hff,8'hfe,8'hf9,8'hf0,8'hf0,8'hf8,8'hfe,8'hfe,8'hfe,8'hfe},
	{8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hf4,8'hf8,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf8,8'hf8,8'hf4,8'hf4,8'hfd},
	{8'hf8,8'hf0,8'hf4,8'hf4,8'hf4,8'hf4,8'hfd,8'hfd,8'hf4,8'hf4,8'hf8,8'hf9,8'hf9,8'hf9,8'hfc,8'hfd,8'hfd,8'hfe,8'hfd,8'hfe,8'hfd,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hfd,8'hf9,8'hf9},
	{8'hfd,8'hf9,8'hf9,8'hf9,8'hf9,8'hfd,8'hf8,8'hf9,8'hfd,8'hf9,8'hfd,8'hfd,8'hf9,8'hfd,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd},
	{8'hf9,8'hfd,8'hfc,8'hfd,8'hf9,8'hfd,8'hf9,8'hf8,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfe,8'hfd,8'hfd,8'hf9},
	{8'hfd,8'hf9,8'hf9,8'hf8,8'hf9,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd},
	{8'hfe,8'hfe,8'hfd,8'hf8,8'hf9,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe},
	{8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe},
	{8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfd,8'hf8,8'hf4,8'hf4,8'hf9,8'hf4,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe},
	{8'h24,8'h24,8'h2d,8'h24,8'h04,8'h00,8'h04,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h25,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h04,8'h04,8'h24},
	{8'h24,8'h00,8'h04,8'h00,8'h24,8'h00,8'h00,8'h25,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24}
	};
	


logic [3:0] wall_type;
//const logic [0:15] [0:15] [3:0] initial_map = '{default:'0}; // for testing purposes

const logic [0:15] [0:15] [3:0]  initial_map = {
 {4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04},
 {4'h04, 4'h02, 4'h02, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h04},
 {4'h04, 4'h02, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h01, 4'h04},
 {4'h04, 4'h00, 4'h00, 4'h04, 4'h00, 4'h00, 4'h04, 4'h00, 4'h00, 4'h04, 4'h00, 4'h00, 4'h04, 4'h00, 4'h01, 4'h04},
 {4'h04, 4'h03, 4'h03, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h02, 4'h00, 4'h00, 4'h00, 4'h00, 4'h04},
 {4'h04, 4'h03, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h02, 4'h00, 4'h00, 4'h00, 4'h00, 4'h04},
 {4'h04, 4'h00, 4'h01, 4'h04, 4'h00, 4'h00, 4'h04, 4'h00, 4'h00, 4'h04, 4'h00, 4'h00, 4'h01, 4'h00, 4'h01, 4'h04},
 {4'h04, 4'h00, 4'h00, 4'h02, 4'h00, 4'h00, 4'h00, 4'h03, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h04},
 {4'h04, 4'h00, 4'h00, 4'h02, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h04},
 {4'h04, 4'h01, 4'h01, 4'h04, 4'h00, 4'h00, 4'h04, 4'h00, 4'h00, 4'h04, 4'h00, 4'h00, 4'h01, 4'h01, 4'h01, 4'h04},
 {4'h04, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h04},
 {4'h04, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h04},
 {4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04, 4'h04},// last line in home screen
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00}};
logic [0:15] [0:15] [3:0]  MazeBitMapMask_p = initial_map;
logic [0:15] [0:15] [3:0]  MazeBitMapMask_n;  

logic [3:0] [0:31][0:31][7:0] object_colors = { wall_4, wall_3, wall_2, wall_1};
 // pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <= TRANSPARENT_ENCODING ;
		MazeBitMapMask_p = initial_map;
		explosion_executed_p <= 0;
	end
	else begin
	explosion_executed_p <= explosion_executed_n;
		RGBout <= TRANSPARENT_ENCODING ; // default 
		MazeBitMapMask_p <= MazeBitMapMask_n;
		if ((InsideRectangle == 1'b1 )		& 	// only if inside the external bracket 
		   (MazeBitMapMask_p[offsetY[8:5] ][offsetX[8:5]] > 4'h0 ))begin
						// take bits 5,6,7,8,9,10 from address to select  position in the maze    
						wall_type = MazeBitMapMask_p[offsetY[8:5] ][offsetX[8:5]] ;
						RGBout <= object_colors[wall_type - 1][offsetY[4:0]][offsetX[4:0]] ; 
		end
	end	
end

always_comb begin 
	increase_score = 0;
	explosion_executed_n = explosion_executed_p;
	MazeBitMapMask_n = MazeBitMapMask_p;
	if (wall_explode && !explosion_executed_p) begin
		if(MazeBitMapMask_p[offsetY[8:5] ][offsetX[8:5]] > 4'h0 && MazeBitMapMask_p[offsetY[8:5] ][offsetX[8:5]] < 4'h4 ) begin
			MazeBitMapMask_n[offsetY[8:5] ][offsetX[8:5]]--; // 
			explosion_executed_n = 1'b1;
			if( MazeBitMapMask_n[offsetY[8:5] ][offsetX[8:5]] == 0 ) // wall destroyed
				increase_score = 1;
		end
	end
	
	if(OneSecPulse) begin
		explosion_executed_n = 0;
	end
	
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule

