// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen Apr  2023  
// (c) Technion IIT, Department of Electrical Engineering 2023 



module	bombMatrixBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic enter_hit, // if enter is hit, put a bomb
					input	 logic signed 	[10:0]	topLeftX, // current position of the player 
					input	 logic signed	[10:0]	topLeftY,  // can be negative , if the object is partliy outside 
					input logic OneSecPulse, 
					input logic addBombCollected,
					
					
					
					output logic [3:0] explosionIndexX,
					output logic [3:0] explosionIndexY,
					output logic explodeBomb,  
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
					
 ) ;
 
 

								 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */


// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 16*16 and use only the top left 16*15 squares 
// this is the bitmap  of the maze , if there is a specific value  the  whole 32*32 rectange will be drawn on the screen
// there are  16 options of differents kinds of 32*32 squares 
// all numbers here are hard coded to simplify the  understanding 


// start the bit map with zeroes, each value represents the timer remaining for the bomb to explode, 0-> no bomb


	const int bomb_timer = 3;
	logic [3:0] max_bomb_limit_p = 3; // number of bombs at the same time
	logic [3:0] max_bomb_limit_n;
   logic [3:0] bomb_counter_p = 0;
	logic [3:0] bomb_counter_n = 0;
	int remaining_time;
	logic bomb_placement_executed_p = 0;
	logic bomb_placement_executed_n = 0;
	
	logic [3:0] explosionIndexX_n;
	logic [3:0] explosionIndexY_n;
	logic explodeBomb_n;
	
	logic [0:15] [0:15] [3:0]  bombBitMapMask_p = '{default:'0}; //don't provide explicit initial values for the array, so it will be initialized with zeroes
	logic [0:15] [0:15] [3:0]  bombBitMapMask_n = '{default:'0};
	// bomb_a is the normal image and bomb_b is a more red version, switching between them gives a dynamic effect.
	const logic [0:31][0:31][7:0] bomb_a = {
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hf9,8'hfc,8'hfc,8'hf8,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hf9,8'he4,8'he0,8'hf8,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hf9,8'hf8,8'hf4,8'hf4,8'hf8,8'hf8,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hf9,8'hf8,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h8d,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h00,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h00,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h00,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h64,8'h64,8'h64,8'hff,8'hff,8'hff,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h00,8'h20,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h20,8'h64,8'h64,8'h64,8'hff,8'hff,8'hff,8'hff,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h24,8'h24,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h64,8'h64,8'h24,8'hff,8'hff,8'hff,8'hff,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h24,8'h24,8'h00,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h00,8'h64,8'h65,8'h24,8'hff,8'hff,8'hff,8'hff,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h24,8'h24,8'h00,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h64,8'h64,8'h64,8'hff,8'hff,8'hff,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h24,8'h24,8'h24,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h64,8'h64,8'h64,8'hff,8'hff,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h24,8'h24,8'h24,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'h00,8'h24,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h24,8'h24,8'h24,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h64,8'h64,8'hff,8'hff,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'h20,8'h00,8'h64,8'hff,8'hff,8'hff,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h24,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h24,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h64,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h00,8'h24,8'h24,8'h24,8'h24,8'h64,8'h64,8'h64,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h20,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff}
	};

 
						
	

	
	
	const logic [0:31][0:31][7:0] bomb_b = {	
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfd,8'hfc,8'hfc,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfd,8'he4,8'he4,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hfd,8'hfc,8'hf8,8'hf8,8'hfc,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'hff,8'hff,8'hff,8'hfd,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'had,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h84,8'h84,8'h84,8'h84,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h20,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h20,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h84,8'h84,8'h84,8'hff,8'hff,8'hff,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h85,8'h20,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h20,8'h84,8'h84,8'h84,8'hff,8'hff,8'hff,8'hff,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h64,8'h64,8'h20,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h84,8'h85,8'h64,8'hff,8'hff,8'hff,8'hff,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h64,8'h64,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h84,8'h8d,8'h64,8'hff,8'hff,8'hff,8'hff,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h64,8'h64,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h84,8'h84,8'h84,8'hff,8'hff,8'hff,8'h85,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h64,8'h64,8'h64,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h84,8'h84,8'h84,8'hff,8'hff,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h64,8'h64,8'h64,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'h20,8'h64,8'h84,8'h84,8'h84,8'h85,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h64,8'h64,8'h64,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h84,8'h84,8'hff,8'hff,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h84,8'hff,8'hff,8'hff,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h64,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h64,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h20,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h84,8'h20,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h84,8'h84,8'h84,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h20,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h64,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff}
	};

	logic[1:0][0:31][0:31][7:0] object_colors = { bomb_b, bomb_a};
	
 
 // pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <= TRANSPARENT_ENCODING ;
		bomb_counter_p <= 0;
	   bombBitMapMask_p <= '{default:'0};
		bomb_placement_executed_p <= 0;
		explodeBomb <= 0;
		explosionIndexX <= 0;
		explosionIndexY <= 0;
		max_bomb_limit_p <= 3;
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 
      bomb_counter_p <= bomb_counter_n;
		bombBitMapMask_p <= bombBitMapMask_n;
		bomb_placement_executed_p <= bomb_placement_executed_n;
		explosionIndexX <= explosionIndexX_n;
		explosionIndexY <= explosionIndexY_n;
		explodeBomb <= explodeBomb_n;
		max_bomb_limit_p <= max_bomb_limit_n;
		remaining_time = bombBitMapMask_p[offsetY[8:5] ][offsetX[8:5]];// take bits 5,6,7,8,9,10 from address to select  position in the maze 
		if ((InsideRectangle == 1'b1 ) && (remaining_time > 4'h00 ))    
						RGBout <= object_colors[remaining_time % 2][offsetY[4:0]][offsetX[4:0]] ; 
		end 
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
always_comb begin

	bomb_counter_n = bomb_counter_p;
	bombBitMapMask_n = bombBitMapMask_p;
	bomb_placement_executed_n = bomb_placement_executed_p;
	explosionIndexX_n = explosionIndexX;
	explosionIndexY_n = explosionIndexY;
	explodeBomb_n = explodeBomb;
	max_bomb_limit_n = max_bomb_limit_p;	
	
	if( (enter_hit == 1'b1) && (bomb_counter_p < max_bomb_limit_p) && (!bomb_placement_executed_p )
		  && (bombBitMapMask_n[topLeftY[8:5] ][topLeftX[8:5]] == 0)	)	begin 	
				bomb_counter_n = bomb_counter_p + 3'b001;
				bombBitMapMask_n[topLeftY[8:5] ][topLeftX[8:5]] = bomb_timer; 
				bomb_placement_executed_n = 1'b1;
	end
	
		if(addBombCollected) begin
			max_bomb_limit_n = 4; // add extra bomb
		end
		
		if ( OneSecPulse ) begin 
			explodeBomb_n = 0;
			bomb_placement_executed_n = 1'b0;
      // Loop through each dimension and initialize to zeroes
			for (int i = 0; i <= 15; i++) begin
				for (int j = 0; j <= 15; j++) begin
						if ( bombBitMapMask_p[i][j] == 4'b0001) begin // bomb about to explode
								bomb_counter_n = bomb_counter_p - 3'b001;
								explosionIndexX_n = j;
								explosionIndexY_n = i;
								explodeBomb_n = 1;
						end 
						if( bombBitMapMask_p[i][j] > 4'b0000) begin
								bombBitMapMask_n[i][j] = bombBitMapMask_p[i][j] - 1; // 1 sec passed, decrement timer 
						end 
				end 
			end 
		end // if OneSecPulse
	
end // start comb
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule

